
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"c1",x"85",x"cb",x"87"),
     1 => (x"ab",x"b7",x"c8",x"83"),
     2 => (x"87",x"c7",x"ff",x"04"),
     3 => (x"26",x"4d",x"26",x"26"),
     4 => (x"26",x"4b",x"26",x"4c"),
     5 => (x"4a",x"71",x"1e",x"4f"),
     6 => (x"5a",x"ce",x"ed",x"c2"),
     7 => (x"48",x"ce",x"ed",x"c2"),
     8 => (x"fe",x"49",x"78",x"c7"),
     9 => (x"4f",x"26",x"87",x"dd"),
    10 => (x"71",x"1e",x"73",x"1e"),
    11 => (x"aa",x"b7",x"c0",x"4a"),
    12 => (x"c2",x"87",x"d3",x"03"),
    13 => (x"05",x"bf",x"f9",x"cd"),
    14 => (x"4b",x"c1",x"87",x"c4"),
    15 => (x"4b",x"c0",x"87",x"c2"),
    16 => (x"5b",x"fd",x"cd",x"c2"),
    17 => (x"cd",x"c2",x"87",x"c4"),
    18 => (x"cd",x"c2",x"5a",x"fd"),
    19 => (x"c1",x"4a",x"bf",x"f9"),
    20 => (x"a2",x"c0",x"c1",x"9a"),
    21 => (x"87",x"e8",x"ec",x"49"),
    22 => (x"cd",x"c2",x"48",x"fc"),
    23 => (x"fe",x"78",x"bf",x"f9"),
    24 => (x"71",x"1e",x"87",x"ef"),
    25 => (x"1e",x"66",x"c4",x"4a"),
    26 => (x"f5",x"e9",x"49",x"72"),
    27 => (x"4f",x"26",x"26",x"87"),
    28 => (x"f9",x"cd",x"c2",x"1e"),
    29 => (x"cf",x"e6",x"49",x"bf"),
    30 => (x"c2",x"ed",x"c2",x"87"),
    31 => (x"78",x"bf",x"e8",x"48"),
    32 => (x"48",x"fe",x"ec",x"c2"),
    33 => (x"c2",x"78",x"bf",x"ec"),
    34 => (x"4a",x"bf",x"c2",x"ed"),
    35 => (x"99",x"ff",x"c3",x"49"),
    36 => (x"72",x"2a",x"b7",x"c8"),
    37 => (x"c2",x"b0",x"71",x"48"),
    38 => (x"26",x"58",x"ca",x"ed"),
    39 => (x"5b",x"5e",x"0e",x"4f"),
    40 => (x"71",x"0e",x"5d",x"5c"),
    41 => (x"87",x"c8",x"ff",x"4b"),
    42 => (x"48",x"fd",x"ec",x"c2"),
    43 => (x"49",x"73",x"50",x"c0"),
    44 => (x"70",x"87",x"f5",x"e5"),
    45 => (x"9c",x"c2",x"4c",x"49"),
    46 => (x"cb",x"49",x"ee",x"cb"),
    47 => (x"49",x"70",x"87",x"c3"),
    48 => (x"fd",x"ec",x"c2",x"4d"),
    49 => (x"c1",x"05",x"bf",x"97"),
    50 => (x"66",x"d0",x"87",x"e2"),
    51 => (x"c6",x"ed",x"c2",x"49"),
    52 => (x"d6",x"05",x"99",x"bf"),
    53 => (x"49",x"66",x"d4",x"87"),
    54 => (x"bf",x"fe",x"ec",x"c2"),
    55 => (x"87",x"cb",x"05",x"99"),
    56 => (x"c3",x"e5",x"49",x"73"),
    57 => (x"02",x"98",x"70",x"87"),
    58 => (x"c1",x"87",x"c1",x"c1"),
    59 => (x"87",x"c0",x"fe",x"4c"),
    60 => (x"d8",x"ca",x"49",x"75"),
    61 => (x"02",x"98",x"70",x"87"),
    62 => (x"ec",x"c2",x"87",x"c6"),
    63 => (x"50",x"c1",x"48",x"fd"),
    64 => (x"97",x"fd",x"ec",x"c2"),
    65 => (x"e3",x"c0",x"05",x"bf"),
    66 => (x"c6",x"ed",x"c2",x"87"),
    67 => (x"66",x"d0",x"49",x"bf"),
    68 => (x"d6",x"ff",x"05",x"99"),
    69 => (x"fe",x"ec",x"c2",x"87"),
    70 => (x"66",x"d4",x"49",x"bf"),
    71 => (x"ca",x"ff",x"05",x"99"),
    72 => (x"e4",x"49",x"73",x"87"),
    73 => (x"98",x"70",x"87",x"c2"),
    74 => (x"87",x"ff",x"fe",x"05"),
    75 => (x"dc",x"fb",x"48",x"74"),
    76 => (x"5b",x"5e",x"0e",x"87"),
    77 => (x"f4",x"0e",x"5d",x"5c"),
    78 => (x"4c",x"4d",x"c0",x"86"),
    79 => (x"c4",x"7e",x"bf",x"ec"),
    80 => (x"ed",x"c2",x"48",x"a6"),
    81 => (x"c1",x"78",x"bf",x"ca"),
    82 => (x"c7",x"1e",x"c0",x"1e"),
    83 => (x"87",x"cd",x"fd",x"49"),
    84 => (x"98",x"70",x"86",x"c8"),
    85 => (x"ff",x"87",x"cd",x"02"),
    86 => (x"87",x"cc",x"fb",x"49"),
    87 => (x"e3",x"49",x"da",x"c1"),
    88 => (x"4d",x"c1",x"87",x"c6"),
    89 => (x"97",x"fd",x"ec",x"c2"),
    90 => (x"87",x"c3",x"02",x"bf"),
    91 => (x"c2",x"87",x"fe",x"d4"),
    92 => (x"4b",x"bf",x"c2",x"ed"),
    93 => (x"bf",x"f9",x"cd",x"c2"),
    94 => (x"87",x"e9",x"c0",x"05"),
    95 => (x"e2",x"49",x"fd",x"c3"),
    96 => (x"fa",x"c3",x"87",x"e6"),
    97 => (x"87",x"e0",x"e2",x"49"),
    98 => (x"ff",x"c3",x"49",x"73"),
    99 => (x"c0",x"1e",x"71",x"99"),
   100 => (x"87",x"ce",x"fb",x"49"),
   101 => (x"b7",x"c8",x"49",x"73"),
   102 => (x"c1",x"1e",x"71",x"29"),
   103 => (x"87",x"c2",x"fb",x"49"),
   104 => (x"fa",x"c5",x"86",x"c8"),
   105 => (x"c6",x"ed",x"c2",x"87"),
   106 => (x"02",x"9b",x"4b",x"bf"),
   107 => (x"cd",x"c2",x"87",x"dd"),
   108 => (x"c7",x"49",x"bf",x"f5"),
   109 => (x"98",x"70",x"87",x"d7"),
   110 => (x"c0",x"87",x"c4",x"05"),
   111 => (x"c2",x"87",x"d2",x"4b"),
   112 => (x"fc",x"c6",x"49",x"e0"),
   113 => (x"f9",x"cd",x"c2",x"87"),
   114 => (x"c2",x"87",x"c6",x"58"),
   115 => (x"c0",x"48",x"f5",x"cd"),
   116 => (x"c2",x"49",x"73",x"78"),
   117 => (x"87",x"cd",x"05",x"99"),
   118 => (x"e1",x"49",x"eb",x"c3"),
   119 => (x"49",x"70",x"87",x"ca"),
   120 => (x"c2",x"02",x"99",x"c2"),
   121 => (x"73",x"4c",x"fb",x"87"),
   122 => (x"05",x"99",x"c1",x"49"),
   123 => (x"f4",x"c3",x"87",x"cd"),
   124 => (x"87",x"f4",x"e0",x"49"),
   125 => (x"99",x"c2",x"49",x"70"),
   126 => (x"fa",x"87",x"c2",x"02"),
   127 => (x"c8",x"49",x"73",x"4c"),
   128 => (x"87",x"cd",x"05",x"99"),
   129 => (x"e0",x"49",x"f5",x"c3"),
   130 => (x"49",x"70",x"87",x"de"),
   131 => (x"d4",x"02",x"99",x"c2"),
   132 => (x"ce",x"ed",x"c2",x"87"),
   133 => (x"87",x"c9",x"02",x"bf"),
   134 => (x"c2",x"88",x"c1",x"48"),
   135 => (x"c2",x"58",x"d2",x"ed"),
   136 => (x"c1",x"4c",x"ff",x"87"),
   137 => (x"c4",x"49",x"73",x"4d"),
   138 => (x"87",x"ce",x"05",x"99"),
   139 => (x"ff",x"49",x"f2",x"c3"),
   140 => (x"70",x"87",x"f5",x"df"),
   141 => (x"02",x"99",x"c2",x"49"),
   142 => (x"ed",x"c2",x"87",x"db"),
   143 => (x"48",x"7e",x"bf",x"ce"),
   144 => (x"03",x"a8",x"b7",x"c7"),
   145 => (x"48",x"6e",x"87",x"cb"),
   146 => (x"ed",x"c2",x"80",x"c1"),
   147 => (x"c2",x"c0",x"58",x"d2"),
   148 => (x"c1",x"4c",x"fe",x"87"),
   149 => (x"49",x"fd",x"c3",x"4d"),
   150 => (x"87",x"cc",x"df",x"ff"),
   151 => (x"99",x"c2",x"49",x"70"),
   152 => (x"c2",x"87",x"d5",x"02"),
   153 => (x"02",x"bf",x"ce",x"ed"),
   154 => (x"c2",x"87",x"c9",x"c0"),
   155 => (x"c0",x"48",x"ce",x"ed"),
   156 => (x"87",x"c2",x"c0",x"78"),
   157 => (x"4d",x"c1",x"4c",x"fd"),
   158 => (x"ff",x"49",x"fa",x"c3"),
   159 => (x"70",x"87",x"e9",x"de"),
   160 => (x"02",x"99",x"c2",x"49"),
   161 => (x"ed",x"c2",x"87",x"d9"),
   162 => (x"c7",x"48",x"bf",x"ce"),
   163 => (x"c0",x"03",x"a8",x"b7"),
   164 => (x"ed",x"c2",x"87",x"c9"),
   165 => (x"78",x"c7",x"48",x"ce"),
   166 => (x"fc",x"87",x"c2",x"c0"),
   167 => (x"c0",x"4d",x"c1",x"4c"),
   168 => (x"c0",x"03",x"ac",x"b7"),
   169 => (x"66",x"c4",x"87",x"d1"),
   170 => (x"82",x"d8",x"c1",x"4a"),
   171 => (x"c6",x"c0",x"02",x"6a"),
   172 => (x"74",x"4b",x"6a",x"87"),
   173 => (x"c0",x"0f",x"73",x"49"),
   174 => (x"1e",x"f0",x"c3",x"1e"),
   175 => (x"f7",x"49",x"da",x"c1"),
   176 => (x"86",x"c8",x"87",x"db"),
   177 => (x"c0",x"02",x"98",x"70"),
   178 => (x"a6",x"c8",x"87",x"e2"),
   179 => (x"ce",x"ed",x"c2",x"48"),
   180 => (x"66",x"c8",x"78",x"bf"),
   181 => (x"c4",x"91",x"cb",x"49"),
   182 => (x"80",x"71",x"48",x"66"),
   183 => (x"bf",x"6e",x"7e",x"70"),
   184 => (x"87",x"c8",x"c0",x"02"),
   185 => (x"c8",x"4b",x"bf",x"6e"),
   186 => (x"0f",x"73",x"49",x"66"),
   187 => (x"c0",x"02",x"9d",x"75"),
   188 => (x"ed",x"c2",x"87",x"c8"),
   189 => (x"f3",x"49",x"bf",x"ce"),
   190 => (x"cd",x"c2",x"87",x"c9"),
   191 => (x"c0",x"02",x"bf",x"fd"),
   192 => (x"c2",x"49",x"87",x"dd"),
   193 => (x"98",x"70",x"87",x"c7"),
   194 => (x"87",x"d3",x"c0",x"02"),
   195 => (x"bf",x"ce",x"ed",x"c2"),
   196 => (x"87",x"ef",x"f2",x"49"),
   197 => (x"cf",x"f4",x"49",x"c0"),
   198 => (x"fd",x"cd",x"c2",x"87"),
   199 => (x"f4",x"78",x"c0",x"48"),
   200 => (x"87",x"e9",x"f3",x"8e"),
   201 => (x"5c",x"5b",x"5e",x"0e"),
   202 => (x"71",x"1e",x"0e",x"5d"),
   203 => (x"ca",x"ed",x"c2",x"4c"),
   204 => (x"cd",x"c1",x"49",x"bf"),
   205 => (x"d1",x"c1",x"4d",x"a1"),
   206 => (x"74",x"7e",x"69",x"81"),
   207 => (x"87",x"cf",x"02",x"9c"),
   208 => (x"74",x"4b",x"a5",x"c4"),
   209 => (x"ca",x"ed",x"c2",x"7b"),
   210 => (x"c8",x"f3",x"49",x"bf"),
   211 => (x"74",x"7b",x"6e",x"87"),
   212 => (x"87",x"c4",x"05",x"9c"),
   213 => (x"87",x"c2",x"4b",x"c0"),
   214 => (x"49",x"73",x"4b",x"c1"),
   215 => (x"d4",x"87",x"c9",x"f3"),
   216 => (x"87",x"c7",x"02",x"66"),
   217 => (x"70",x"87",x"da",x"49"),
   218 => (x"c0",x"87",x"c2",x"4a"),
   219 => (x"c1",x"ce",x"c2",x"4a"),
   220 => (x"d8",x"f2",x"26",x"5a"),
   221 => (x"00",x"00",x"00",x"87"),
   222 => (x"00",x"00",x"00",x"00"),
   223 => (x"00",x"00",x"00",x"00"),
   224 => (x"4a",x"71",x"1e",x"00"),
   225 => (x"49",x"bf",x"c8",x"ff"),
   226 => (x"26",x"48",x"a1",x"72"),
   227 => (x"c8",x"ff",x"1e",x"4f"),
   228 => (x"c0",x"fe",x"89",x"bf"),
   229 => (x"c0",x"c0",x"c0",x"c0"),
   230 => (x"87",x"c4",x"01",x"a9"),
   231 => (x"87",x"c2",x"4a",x"c0"),
   232 => (x"48",x"72",x"4a",x"c1"),
   233 => (x"5e",x"0e",x"4f",x"26"),
   234 => (x"0e",x"5d",x"5c",x"5b"),
   235 => (x"d4",x"ff",x"4b",x"71"),
   236 => (x"48",x"66",x"d0",x"4c"),
   237 => (x"49",x"d6",x"78",x"c0"),
   238 => (x"87",x"ec",x"db",x"ff"),
   239 => (x"6c",x"7c",x"ff",x"c3"),
   240 => (x"99",x"ff",x"c3",x"49"),
   241 => (x"c3",x"49",x"4d",x"71"),
   242 => (x"e0",x"c1",x"99",x"f0"),
   243 => (x"87",x"cb",x"05",x"a9"),
   244 => (x"6c",x"7c",x"ff",x"c3"),
   245 => (x"d0",x"98",x"c3",x"48"),
   246 => (x"c3",x"78",x"08",x"66"),
   247 => (x"4a",x"6c",x"7c",x"ff"),
   248 => (x"c3",x"31",x"c8",x"49"),
   249 => (x"4a",x"6c",x"7c",x"ff"),
   250 => (x"49",x"72",x"b2",x"71"),
   251 => (x"ff",x"c3",x"31",x"c8"),
   252 => (x"71",x"4a",x"6c",x"7c"),
   253 => (x"c8",x"49",x"72",x"b2"),
   254 => (x"7c",x"ff",x"c3",x"31"),
   255 => (x"b2",x"71",x"4a",x"6c"),
   256 => (x"c0",x"48",x"d0",x"ff"),
   257 => (x"9b",x"73",x"78",x"e0"),
   258 => (x"72",x"87",x"c2",x"02"),
   259 => (x"26",x"48",x"75",x"7b"),
   260 => (x"26",x"4c",x"26",x"4d"),
   261 => (x"1e",x"4f",x"26",x"4b"),
   262 => (x"5e",x"0e",x"4f",x"26"),
   263 => (x"f8",x"0e",x"5c",x"5b"),
   264 => (x"c8",x"1e",x"76",x"86"),
   265 => (x"fd",x"fd",x"49",x"a6"),
   266 => (x"70",x"86",x"c4",x"87"),
   267 => (x"c8",x"48",x"6e",x"4b"),
   268 => (x"c6",x"c3",x"03",x"a8"),
   269 => (x"c3",x"4a",x"73",x"87"),
   270 => (x"d0",x"c1",x"9a",x"f0"),
   271 => (x"87",x"c7",x"02",x"aa"),
   272 => (x"05",x"aa",x"e0",x"c1"),
   273 => (x"73",x"87",x"f4",x"c2"),
   274 => (x"02",x"99",x"c8",x"49"),
   275 => (x"c6",x"ff",x"87",x"c3"),
   276 => (x"c3",x"4c",x"73",x"87"),
   277 => (x"05",x"ac",x"c2",x"9c"),
   278 => (x"c4",x"87",x"cd",x"c1"),
   279 => (x"31",x"c9",x"49",x"66"),
   280 => (x"66",x"c4",x"1e",x"71"),
   281 => (x"c2",x"92",x"d4",x"4a"),
   282 => (x"72",x"49",x"d2",x"ed"),
   283 => (x"fe",x"d4",x"fe",x"81"),
   284 => (x"49",x"66",x"c4",x"87"),
   285 => (x"49",x"e3",x"c0",x"1e"),
   286 => (x"87",x"d1",x"d9",x"ff"),
   287 => (x"d8",x"ff",x"49",x"d8"),
   288 => (x"c0",x"c8",x"87",x"e6"),
   289 => (x"c2",x"dc",x"c2",x"1e"),
   290 => (x"ce",x"f1",x"fd",x"49"),
   291 => (x"48",x"d0",x"ff",x"87"),
   292 => (x"c2",x"78",x"e0",x"c0"),
   293 => (x"d0",x"1e",x"c2",x"dc"),
   294 => (x"92",x"d4",x"4a",x"66"),
   295 => (x"49",x"d2",x"ed",x"c2"),
   296 => (x"d3",x"fe",x"81",x"72"),
   297 => (x"86",x"d0",x"87",x"c6"),
   298 => (x"c1",x"05",x"ac",x"c1"),
   299 => (x"66",x"c4",x"87",x"cd"),
   300 => (x"71",x"31",x"c9",x"49"),
   301 => (x"4a",x"66",x"c4",x"1e"),
   302 => (x"ed",x"c2",x"92",x"d4"),
   303 => (x"81",x"72",x"49",x"d2"),
   304 => (x"87",x"eb",x"d3",x"fe"),
   305 => (x"1e",x"c2",x"dc",x"c2"),
   306 => (x"d4",x"4a",x"66",x"c8"),
   307 => (x"d2",x"ed",x"c2",x"92"),
   308 => (x"fe",x"81",x"72",x"49"),
   309 => (x"c8",x"87",x"d2",x"d1"),
   310 => (x"c0",x"1e",x"49",x"66"),
   311 => (x"d7",x"ff",x"49",x"e3"),
   312 => (x"49",x"d7",x"87",x"eb"),
   313 => (x"87",x"c0",x"d7",x"ff"),
   314 => (x"c2",x"1e",x"c0",x"c8"),
   315 => (x"fd",x"49",x"c2",x"dc"),
   316 => (x"d0",x"87",x"d2",x"ef"),
   317 => (x"48",x"d0",x"ff",x"86"),
   318 => (x"f8",x"78",x"e0",x"c0"),
   319 => (x"87",x"d1",x"fc",x"8e"),
   320 => (x"5c",x"5b",x"5e",x"0e"),
   321 => (x"71",x"1e",x"0e",x"5d"),
   322 => (x"4c",x"d4",x"ff",x"4d"),
   323 => (x"48",x"7e",x"66",x"d4"),
   324 => (x"06",x"a8",x"b7",x"c3"),
   325 => (x"48",x"c0",x"87",x"c5"),
   326 => (x"75",x"87",x"e2",x"c1"),
   327 => (x"df",x"e1",x"fe",x"49"),
   328 => (x"c4",x"1e",x"75",x"87"),
   329 => (x"93",x"d4",x"4b",x"66"),
   330 => (x"83",x"d2",x"ed",x"c2"),
   331 => (x"cc",x"fe",x"49",x"73"),
   332 => (x"83",x"c8",x"87",x"db"),
   333 => (x"d0",x"ff",x"4b",x"6b"),
   334 => (x"78",x"e1",x"c8",x"48"),
   335 => (x"49",x"73",x"7c",x"dd"),
   336 => (x"71",x"99",x"ff",x"c3"),
   337 => (x"c8",x"49",x"73",x"7c"),
   338 => (x"ff",x"c3",x"29",x"b7"),
   339 => (x"73",x"7c",x"71",x"99"),
   340 => (x"29",x"b7",x"d0",x"49"),
   341 => (x"71",x"99",x"ff",x"c3"),
   342 => (x"d8",x"49",x"73",x"7c"),
   343 => (x"7c",x"71",x"29",x"b7"),
   344 => (x"7c",x"7c",x"7c",x"c0"),
   345 => (x"7c",x"7c",x"7c",x"7c"),
   346 => (x"7c",x"7c",x"7c",x"7c"),
   347 => (x"78",x"e0",x"c0",x"7c"),
   348 => (x"dc",x"1e",x"66",x"c4"),
   349 => (x"d4",x"d5",x"ff",x"49"),
   350 => (x"73",x"86",x"c8",x"87"),
   351 => (x"ce",x"fa",x"26",x"48"),
   352 => (x"5b",x"5e",x"0e",x"87"),
   353 => (x"1e",x"0e",x"5d",x"5c"),
   354 => (x"d4",x"ff",x"7e",x"71"),
   355 => (x"c2",x"1e",x"6e",x"4b"),
   356 => (x"fe",x"49",x"f2",x"ef"),
   357 => (x"c4",x"87",x"f6",x"ca"),
   358 => (x"9d",x"4d",x"70",x"86"),
   359 => (x"87",x"c3",x"c3",x"02"),
   360 => (x"bf",x"fa",x"ef",x"c2"),
   361 => (x"fe",x"49",x"6e",x"4c"),
   362 => (x"ff",x"87",x"d5",x"df"),
   363 => (x"c5",x"c8",x"48",x"d0"),
   364 => (x"7b",x"d6",x"c1",x"78"),
   365 => (x"7b",x"15",x"4a",x"c0"),
   366 => (x"e0",x"c0",x"82",x"c1"),
   367 => (x"f5",x"04",x"aa",x"b7"),
   368 => (x"48",x"d0",x"ff",x"87"),
   369 => (x"c5",x"c8",x"78",x"c4"),
   370 => (x"7b",x"d3",x"c1",x"78"),
   371 => (x"78",x"c4",x"7b",x"c1"),
   372 => (x"c1",x"02",x"9c",x"74"),
   373 => (x"dc",x"c2",x"87",x"fc"),
   374 => (x"c0",x"c8",x"7e",x"c2"),
   375 => (x"b7",x"c0",x"8c",x"4d"),
   376 => (x"87",x"c6",x"03",x"ac"),
   377 => (x"4d",x"a4",x"c0",x"c8"),
   378 => (x"e8",x"c2",x"4c",x"c0"),
   379 => (x"49",x"bf",x"97",x"f3"),
   380 => (x"d2",x"02",x"99",x"d0"),
   381 => (x"c2",x"1e",x"c0",x"87"),
   382 => (x"fe",x"49",x"f2",x"ef"),
   383 => (x"c4",x"87",x"ea",x"cc"),
   384 => (x"4a",x"49",x"70",x"86"),
   385 => (x"c2",x"87",x"ef",x"c0"),
   386 => (x"c2",x"1e",x"c2",x"dc"),
   387 => (x"fe",x"49",x"f2",x"ef"),
   388 => (x"c4",x"87",x"d6",x"cc"),
   389 => (x"4a",x"49",x"70",x"86"),
   390 => (x"c8",x"48",x"d0",x"ff"),
   391 => (x"d4",x"c1",x"78",x"c5"),
   392 => (x"bf",x"97",x"6e",x"7b"),
   393 => (x"c1",x"48",x"6e",x"7b"),
   394 => (x"c1",x"7e",x"70",x"80"),
   395 => (x"f0",x"ff",x"05",x"8d"),
   396 => (x"48",x"d0",x"ff",x"87"),
   397 => (x"9a",x"72",x"78",x"c4"),
   398 => (x"c0",x"87",x"c5",x"05"),
   399 => (x"87",x"e5",x"c0",x"48"),
   400 => (x"ef",x"c2",x"1e",x"c1"),
   401 => (x"c9",x"fe",x"49",x"f2"),
   402 => (x"86",x"c4",x"87",x"fe"),
   403 => (x"fe",x"05",x"9c",x"74"),
   404 => (x"d0",x"ff",x"87",x"c4"),
   405 => (x"78",x"c5",x"c8",x"48"),
   406 => (x"c0",x"7b",x"d3",x"c1"),
   407 => (x"c1",x"78",x"c4",x"7b"),
   408 => (x"c0",x"87",x"c2",x"48"),
   409 => (x"4d",x"26",x"26",x"48"),
   410 => (x"4b",x"26",x"4c",x"26"),
   411 => (x"5e",x"0e",x"4f",x"26"),
   412 => (x"71",x"0e",x"5c",x"5b"),
   413 => (x"02",x"66",x"cc",x"4b"),
   414 => (x"c0",x"4c",x"87",x"d8"),
   415 => (x"d8",x"02",x"8c",x"f0"),
   416 => (x"c1",x"4a",x"74",x"87"),
   417 => (x"87",x"d1",x"02",x"8a"),
   418 => (x"87",x"cd",x"02",x"8a"),
   419 => (x"87",x"c9",x"02",x"8a"),
   420 => (x"49",x"73",x"87",x"d7"),
   421 => (x"d0",x"87",x"ea",x"fb"),
   422 => (x"c0",x"1e",x"74",x"87"),
   423 => (x"87",x"e0",x"f9",x"49"),
   424 => (x"49",x"73",x"1e",x"74"),
   425 => (x"c8",x"87",x"d9",x"f9"),
   426 => (x"87",x"fc",x"fe",x"86"),
   427 => (x"db",x"c2",x"1e",x"00"),
   428 => (x"c1",x"49",x"bf",x"d6"),
   429 => (x"da",x"db",x"c2",x"b9"),
   430 => (x"48",x"d4",x"ff",x"59"),
   431 => (x"ff",x"78",x"ff",x"c3"),
   432 => (x"e1",x"c8",x"48",x"d0"),
   433 => (x"48",x"d4",x"ff",x"78"),
   434 => (x"31",x"c4",x"78",x"c1"),
   435 => (x"d0",x"ff",x"78",x"71"),
   436 => (x"78",x"e0",x"c0",x"48"),
   437 => (x"00",x"00",x"4f",x"26"),
   438 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

